module sreg4 {
    
}